// ========================================================================================
//
// File:             multiplier.sv
// Description:      A 32-bit signed multiplier module
// Author:           Aaron Pitcher (pitchea@mcmaster.ca)
// Date:             07-Jun-2021 03:18:11 PM
//
// Copyright 2021 Aaron Pitcher
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//
// ========================================================================================
`timescale 1ns/100ps

module multiplier #(
    parameter WIDTH = 32
)(
    input logic [WIDTH-1:0] op1,
    input logic [WIDTH-1:0] op2,
    output logic [WIDTH-1:0] result
);

    logic [2*WIDTH-1:0] result_long;

    assign result_long = $signed(op1) * $signed(op2);
    assign result = result_long[WIDTH-1:0];

endmodule

// ========================================================================================
// EoF
// ========================================================================================